//////////////////////////////////////
//  Author: YiBo Zhang
//  Date: 2022-03-14 14:09:50
//  LastEditTime: 2022-03-14 14:15:15
//  LastEditors: YiBo Zhang
//  Description: this is alu
//  
 /////////////////////////////////////
module fb_alu (
  input [1:0] alu_op,
  input [`FB_32BITS-1:0] op1,
  input [`FB_32BITS-1:0] op2,
  output [`FB_32BITS-1:0] alu_res
);
  
endmodule