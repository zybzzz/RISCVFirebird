// `include "../../rtl/fb_regfile.v"
module tb_test;

initial begin
  $display("hello world!");
  $finish;
end

endmodule
